module LSB_Four_AproximateORAdder(
  input [7:0] A,
  input [7:0] B,
  input Cin,
  output [7:0] S,
  output Cout);

wire cin, cout1,cout2,cout3, cout4, cout5, cout6, cout7;

assign S[7] = A[7] | B[7];
assign S[6] = A[6] | B[6];
assign S[5] = A[5] | B[5];
assign S[4] = A[4] | B[4];
assign cin = A[4] & B[4];
FullAdder fa3 (A[3], B[3], cin, S[3], cout3);
FullAdder fa2 (A[2], B[2], cout3, S[2], cout2);
FullAdder fa1 (A[1], B[1], cout2, S[1], cout1);
FullAdder fa0 (A[0], B[0], cout1, S[0], Cout);

endmodule
